module io(input [15:0] io_dip, output [15:0] io_led);
    assign io_led = io_dip;
endmodule