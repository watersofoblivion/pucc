/*
 * A UART Receiver
 */