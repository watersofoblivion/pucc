/*
 * A UART Transmitter
 */