/*
 * A UART
 */