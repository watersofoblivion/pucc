/**
 */
module HDubCoreLogicAny#(WIDTH = 1)(HDubCoreLogicUnOpIf.Impl iface);
endmodule
