interface Shifter;
endinterface;

/*
 * Implementation
 */

module ShifterImpl(Shifter.Impl iface, ShiftLeftLogical.Injected sll, ShiftRightLogical.Injected srl, ShiftRightArithmetic.Injected sra);
endmodule;