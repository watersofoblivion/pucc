module HDubCoreLogicAll#(WIDTH = 1)(HDubCoreLogicUnOpIf.Impl iface);
endmodule
