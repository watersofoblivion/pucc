module HDubCoreLogicBitwiseAndOp #(WIDTH = 1);
endmodule
