module HDubCoreLogicBitwiseOrOp #(WIDTH = 1);
endmodule
