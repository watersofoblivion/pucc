module HDubCoreLogicBitwiseNotOp #(WIDTH = 1);
endmodule