module HDubCoreLogicBitwiseXorOp #(WIDTH = 1);
endmodule
