package hdub_core_logic_gate;
    typedef enum {
        GATE_AND,
        GATE_OR,
        GATE_NOT,
        GATE_XOR
    } gate_type;
endpackage
