/*
 * A FIFO
 */