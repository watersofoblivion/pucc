module HDubCoreLogicNone#(WIDTH = 1)(HDubCoreLogicUnOpIf.Impl iface);
endmodule
